`ifndef COMMON_DEFINES_SVH
`define COMMON_DEFINES_SVH

`define DATA_WIDTH 64
`define INSTR_WIDTH 32
`define RAM_REAL_SIZE 10

`define REG_ADDR_WIDTH 5

`endif